`default_nettype none

module task2_fsm(clk, s, done_flag);
endmodule