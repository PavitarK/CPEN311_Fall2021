module swap_fsm(clk, counter_i, counter_j, s);
endmodule